*.include "/home/ff/eecs251b/sky130/sky130_cds/sky130_release_0.0.1/models/sky130.lib.spice" section=tt
*.include "/home/ff/eecs251b/sky130/sky130_cds/sky130_release_0.0.1/models/sky130.lib.spice" tt
*.include '/home/ff/eecs251b/sky130/sky130_conv.spice'

.SUBCKT coarse_pass_transistors Vgn_0 Vgn_1 Vgn_2 Vgn_3 Vgn_4 Vgn_5 Vgn_6 Vgn_7 Vgn_8 Vgn_9 Vgn_10 Vgn_11 Vgn_12 Vgn_13 Vgn_14 Vgn_15 Vout VDD VSS
   
   Xinst257 Vgn_0 VSS VSS VDD VDD Vg_0 sky130_fd_sc_hd__inv_16
   Xinst258 Vgn_1 VSS VSS VDD VDD Vg_1 sky130_fd_sc_hd__inv_16
   Xinst259 Vgn_2 VSS VSS VDD VDD Vg_2 sky130_fd_sc_hd__inv_16
   Xinst260 Vgn_3 VSS VSS VDD VDD Vg_3 sky130_fd_sc_hd__inv_16
   Xinst261 Vgn_4 VSS VSS VDD VDD Vg_4 sky130_fd_sc_hd__inv_16
   Xinst262 Vgn_5 VSS VSS VDD VDD Vg_5 sky130_fd_sc_hd__inv_16 
   Xinst263 Vgn_6 VSS VSS VDD VDD Vg_6 sky130_fd_sc_hd__inv_16
   Xinst264 Vgn_7 VSS VSS VDD VDD Vg_7 sky130_fd_sc_hd__inv_16 
   Xinst265 Vgn_8 VSS VSS VDD VDD Vg_8 sky130_fd_sc_hd__inv_16
   Xinst266 Vgn_9 VSS VSS VDD VDD Vg_9 sky130_fd_sc_hd__inv_16
   Xinst267 Vgn_10 VSS VSS VDD VDD Vg_10 sky130_fd_sc_hd__inv_16
   Xinst268 Vgn_11 VSS VSS VDD VDD Vg_11 sky130_fd_sc_hd__inv_16
   Xinst269 Vgn_12 VSS VSS VDD VDD Vg_12 sky130_fd_sc_hd__inv_16
   Xinst270 Vgn_13 VSS VSS VDD VDD Vg_13 sky130_fd_sc_hd__inv_16 
   Xinst271 Vgn_14 VSS VSS VDD VDD Vg_14 sky130_fd_sc_hd__inv_16
   Xinst272 Vgn_15 VSS VSS VDD VDD Vg_15 sky130_fd_sc_hd__inv_16 
   Xinst1 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst2 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst3 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst4 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst5 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst6 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst7 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst8 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst9 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst10 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst11 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst12 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst13 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst14 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst15 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst16 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u

   Xinst17 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst18 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst19 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst20 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst21 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst22 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst23 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst24 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst25 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst26 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst27 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst28 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst29 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst30 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst31 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst32 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u

   Xinst33 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst34 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst35 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst36 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst37 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst38 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst39 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst40 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst41 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst42 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst43 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst44 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst45 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst46 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst47 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst48 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst49 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst50 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst51 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst52 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst53 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst54 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst55 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst56 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst57 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst58 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst59 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst60 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst61 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst62 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst63 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst64 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst65 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst66 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst67 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst68 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst69 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst70 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst71 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst72 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst73 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst74 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst75 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst76 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst77 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst78 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst79 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst80 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst81 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst82 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst83 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst84 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst85 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst86 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst87 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst88 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst89 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst90 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst91 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst92 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst93 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst94 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst95 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst96 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst97 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst98 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst99 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst100 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst101 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst102 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst103 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst104 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst105 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst106 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst107 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst108 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst109 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst110 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst111 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst112 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst113 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst114 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst115 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst116 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst117 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst118 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst119 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst120 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst121 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst122 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst123 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst124 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst125 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst126 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst127 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst128 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst129 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst130 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst131 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst132 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst133 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst134 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst135 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst136 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst137 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst138 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst139 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst140 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst141 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst142 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst143 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst144 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst145 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst146 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst147 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst148 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst149 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst150 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst151 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst152 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst153 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst154 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst155 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst156 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst157 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst158 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst159 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst160 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst161 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst162 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst163 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst164 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst165 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst166 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst167 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst168 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst169 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst170 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst171 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst172 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst173 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst174 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst175 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst176 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst177 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst178 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst179 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst180 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst181 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst182 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst183 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst184 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst185 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst186 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst187 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst188 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst189 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst190 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst191 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst192 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst193 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst194 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst195 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst196 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst197 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst198 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst199 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst200 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst201 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst202 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst203 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst204 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst205 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst206 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst207 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst208 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst209 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst210 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst211 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst212 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst213 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst214 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst215 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst216 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst217 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst218 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst219 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst220 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst221 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst222 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst223 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst224 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst225 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst226 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst227 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst228 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst229 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst230 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst231 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst232 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst233 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst234 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst235 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst236 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst237 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst238 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst239 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst240 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
   Xinst241 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst242 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst243 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst244 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst245 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst246 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst247 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst248 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst249 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst250 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst251 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst252 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst253 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst254 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst255 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst256 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u

.ENDS coarse_pass_transistors
