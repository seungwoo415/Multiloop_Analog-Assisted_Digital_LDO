
.SUBCKT pass_transistors_256 vg0 vg1 vg2 vg3 vg4 vg5 vg6 vg7 vg8 vg9 vg10 vg11 vg12 vg13 vg14 vg15 vg16 vg17 vg18 vg19 vg20 vg21 vg22 vg23 vg24 vg25 vg26 vg27 vg28 vg29 vg30 vg31 vg32 vg33 vg34 vg35 vg36 vg37 vg38 vg39 vg40 vg41 vg42 vg43 vg44 vg45 vg46 vg47 vg48 vg49 vg50 vg51 vg52 vg53 vg54 vg55 vg56 vg57 vg58 vg59 vg60 vg61 vg62 vg63 vg64 vg65 vg66 vg67 vg68 vg69 vg70 vg71 vg72 vg73 vg74 vg75 vg76 vg77 vg78 vg79 vg80 vg81 vg82 vg83 vg84 vg85 vg86 vg87 vg88 vg89 vg90 vg91 vg92 vg93 vg94 vg95 vg96 vg97 vg98 vg99 vg100 vg101 vg102 vg103 vg104 vg105 vg106 vg107 vg108 vg109 vg110 vg111 vg112 vg113 vg114 vg115 vg116 vg117 vg118 vg119 vg120 vg121 vg122 vg123 vg124 vg125 vg126 vg127 vg128 vg129 vg130 vg131 vg132 vg133 vg134 vg135 vg136 vg137 vg138 vg139 vg140 vg141 vg142 vg143 vg144 vg145 vg146 vg147 vg148 vg149 vg150 vg151 vg152 vg153 vg154 vg155 vg156 vg157 vg158 vg159 vg160 vg161 vg162 vg163 vg164 vg165 vg166 vg167 vg168 vg169 vg170 vg171 vg172 vg173 vg174 vg175 vg176 vg177 vg178 vg179 vg180 vg181 vg182 vg183 vg184 vg185 vg186 vg187 vg188 vg189 vg190 vg191 vg192 vg193 vg194 vg195 vg196 vg197 vg198 vg199 vg200 vg201 vg202 vg203 vg204 vg205 vg206 vg207 vg208 vg209 vg210 vg211 vg212 vg213 vg214 vg215 vg216 vg217 vg218 vg219 vg220 vg221 vg222 vg223 vg224 vg225 vg226 vg227 vg228 vg229 vg230 vg231 vg232 vg233 vg234 vg235 vg236 vg237 vg238 vg239 vg240 vg241 vg242 vg243 vg244 vg245 vg246 vg247 vg248 vg249 vg250 vg251 vg252 vg253 vg254 vg255 vout vdd 
 
   Xinst1 vout vg0 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst2 vout vg1 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst3 vout vg2 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst4 vout vg3 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst5 vout vg4 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst6 vout vg5 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst7 vout vg6 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst8 vout vg7 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst9 vout vg8 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst10 vout vg9 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst11 vout vg10 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst12 vout vg11 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst13 vout vg12 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst14 vout vg13 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst15 vout vg14 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst16 vout vg15 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst17 vout vg16 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst18 vout vg17 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst19 vout vg18 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst20 vout vg19 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst21 vout vg20 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst22 vout vg21 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst23 vout vg22 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst24 vout vg23 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst25 vout vg24 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst26 vout vg25 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst27 vout vg26 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst28 vout vg27 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst29 vout vg28 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst30 vout vg29 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst31 vout vg30 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst32 vout vg31 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst33 vout vg32 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst34 vout vg33 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst35 vout vg34 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst36 vout vg35 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst37 vout vg36 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst38 vout vg37 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst39 vout vg38 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst40 vout vg39 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst41 vout vg40 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst42 vout vg41 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst43 vout vg42 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst44 vout vg43 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst45 vout vg44 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst46 vout vg45 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst47 vout vg46 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst48 vout vg47 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst49 vout vg48 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst50 vout vg49 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst51 vout vg50 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst52 vout vg51 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst53 vout vg52 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst54 vout vg53 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst55 vout vg54 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst56 vout vg55 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst57 vout vg56 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst58 vout vg57 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst59 vout vg58 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst60 vout vg59 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst61 vout vg60 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst62 vout vg61 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst63 vout vg62 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst64 vout vg63 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst65 vout vg64 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst66 vout vg65 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst67 vout vg66 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst68 vout vg67 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst69 vout vg68 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst70 vout vg69 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst71 vout vg70 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst72 vout vg71 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst73 vout vg72 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst74 vout vg73 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst75 vout vg74 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst76 vout vg75 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst77 vout vg76 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst78 vout vg77 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst79 vout vg78 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst80 vout vg79 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst81 vout vg80 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst82 vout vg81 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst83 vout vg82 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst84 vout vg83 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst85 vout vg84 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst86 vout vg85 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst87 vout vg86 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst88 vout vg87 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst89 vout vg88 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst90 vout vg89 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst91 vout vg90 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst92 vout vg91 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst93 vout vg92 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst94 vout vg93 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst95 vout vg94 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst96 vout vg95 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst97 vout vg96 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst98 vout vg97 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst99 vout vg98 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst100 vout vg99 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst101 vout vg100 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst102 vout vg101 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst103 vout vg102 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst104 vout vg103 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst105 vout vg104 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst106 vout vg105 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst107 vout vg106 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst108 vout vg107 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst109 vout vg108 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst110 vout vg109 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst111 vout vg110 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst112 vout vg111 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst113 vout vg112 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst114 vout vg113 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst115 vout vg114 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst116 vout vg115 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst117 vout vg116 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst118 vout vg117 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst119 vout vg118 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst120 vout vg119 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst121 vout vg120 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst122 vout vg121 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst123 vout vg122 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst124 vout vg123 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst125 vout vg124 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst126 vout vg125 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst127 vout vg126 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst128 vout vg127 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst129 vout vg128 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst130 vout vg129 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst131 vout vg130 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst132 vout vg131 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst133 vout vg132 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst134 vout vg133 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst135 vout vg134 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst136 vout vg135 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst137 vout vg136 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst138 vout vg137 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst139 vout vg138 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst140 vout vg139 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst141 vout vg140 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst142 vout vg141 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst143 vout vg142 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst144 vout vg143 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst145 vout vg144 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst146 vout vg145 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst147 vout vg146 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst148 vout vg147 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst149 vout vg148 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst150 vout vg149 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst151 vout vg150 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst152 vout vg151 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst153 vout vg152 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst154 vout vg153 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst155 vout vg154 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst156 vout vg155 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst157 vout vg156 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst158 vout vg157 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst159 vout vg158 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst160 vout vg159 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst161 vout vg160 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst162 vout vg161 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst163 vout vg162 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst164 vout vg163 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst165 vout vg164 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst166 vout vg165 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst167 vout vg166 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst168 vout vg167 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst169 vout vg168 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst170 vout vg169 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst171 vout vg170 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst172 vout vg171 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst173 vout vg172 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst174 vout vg173 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst175 vout vg174 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst176 vout vg175 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst177 vout vg176 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst178 vout vg177 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst179 vout vg178 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst180 vout vg179 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst181 vout vg180 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst182 vout vg181 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst183 vout vg182 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst184 vout vg183 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst185 vout vg184 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst186 vout vg185 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst187 vout vg186 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst188 vout vg187 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst189 vout vg188 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst190 vout vg189 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst191 vout vg190 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst192 vout vg191 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst193 vout vg192 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst194 vout vg193 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst195 vout vg194 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst196 vout vg195 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst197 vout vg196 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst198 vout vg197 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst199 vout vg198 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst200 vout vg199 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst201 vout vg200 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst202 vout vg201 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst203 vout vg202 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst204 vout vg203 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst205 vout vg204 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst206 vout vg205 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst207 vout vg206 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst208 vout vg207 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst209 vout vg208 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst210 vout vg209 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst211 vout vg210 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst212 vout vg211 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst213 vout vg212 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst214 vout vg213 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst215 vout vg214 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst216 vout vg215 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst217 vout vg216 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst218 vout vg217 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst219 vout vg218 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst220 vout vg219 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst221 vout vg220 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst222 vout vg221 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst223 vout vg222 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst224 vout vg223 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst225 vout vg224 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst226 vout vg225 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst227 vout vg226 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst228 vout vg227 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst229 vout vg228 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst230 vout vg229 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst231 vout vg230 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst232 vout vg231 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst233 vout vg232 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst234 vout vg233 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst235 vout vg234 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst236 vout vg235 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst237 vout vg236 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst238 vout vg237 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst239 vout vg238 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst240 vout vg239 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst241 vout vg240 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst242 vout vg241 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst243 vout vg242 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst244 vout vg243 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst245 vout vg244 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst246 vout vg245 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst247 vout vg246 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst248 vout vg247 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst249 vout vg248 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst250 vout vg249 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst251 vout vg250 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst252 vout vg251 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst253 vout vg252 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst254 vout vg253 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst255 vout vg254 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   Xinst256 vout vg255 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=0.5u
   
.ENDS pass_transistors_256
