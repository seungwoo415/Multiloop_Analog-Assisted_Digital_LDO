
.include './../strong_arm_system.sp'
.include 'dllogic.sp' 
.include 'pass_transistors_256.sp'  
*.include '/home/aa/users/cs199-apt/Downloads/sky130_fd_sc_hd.spice' 
*.include '/home/ff/eecs251b/sky130/sky130_cds/sky130_release_0.0.1/models/sky130.lib.spice'
*.include '/home/ff/eecs251b/sky130/sky130_conv.spice'

.SUBCKT ldo_core ldotop_vref ldotop_vdd ldotop_vss ldotop_clk ldotop_rst ldotop_vout  

  xinst0 ldotop_vref ldotop_vout output_p output_n real_clk ldotop_vdd ldotop_vss strong_arm_system
  xinst5 ldotop_vdd ldotop_vss ldotop_clk real_clk inverter 
  xinst1 ldotop_vdd ldotop_vss output_p real_output inverter
  xinst2 ldotop_vdd ldotop_vss output_n fake_output inverter
  xinst3 ldotop_clk ldotop_rst fake_output out255 out254 out253 out252 out251 out250 out249 out248 out247 out246 out245 out244 out243 out242 out241 out240 out239 out238 out237 out236 out235 out234 out233 out232 out231 out230 out229 out228 out227 out226 out225 out224 out223 out222 out221 out220 out219 out218 out217 out216 out215 out214 out213 out212 out211 out210 out209 out208 out207 out206 out205 out204 out203 out202 out201 out200 out199 out198 out197 out196 out195 out194 out193 out192 out191 out190 out189 out188 out187 out186 out185 out184 out183 out182 out181 out180 out179 out178 out177 out176 out175 out174 out173 out172 out171 out170 out169 out168 out167 out166 out165 out164 out163 out162 out161 out160 out159 out158 out157 out156 out155 out154 out153 out152 out151 out150 out149 out148 out147 out146 out145 out144 out143 out142 out141 out140 out139 out138 out137 out136 out135 out134 out133 out132 out131 out130 out129 out128 out127 out126 out125 out124 out123 out122 out121 out120 out119 out118 out117 out116 out115 out114 out113 out112 out111 out110 out109 out108 out107 out106 out105 out104 out103 out102 out101 out100 out99 out98 out97 out96 out95 out94 out93 out92 out91 out90 out89 out88 out87 out86 out85 out84 out83 out82 out81 out80 out79 out78 out77 out76 out75 out74 out73 out72 out71 out70 out69 out68 out67 out66 out65 out64 out63 out62 out61 out60 out59 out58 out57 out56 out55 out54 out53 out52 out51 out50 out49 out48 out47 out46 out45 out44 out43 out42 out41 out40 out39 out38 out37 out36 out35 out34 out33 out32 out31 out30 out29 out28 out27 out26 out25 out24 out23 out22 out21 out20 out19 out18 out17 out16 out15 out14 out13 out12 out11 out10 out9 out8 out7 out6 out5 out4 out3 out2 out1 out0 ldotop_vdd ldotop_vss DigitalLDOLogic 
  xinst4 out255 out254 out253 out252 out251 out250 out249 out248 out247 out246 out245 out244 out243 out242 out241 out240 out239 out238 out237 out236 out235 out234 out233 out232 out231 out230 out229 out228 out227 out226 out225 out224 out223 out222 out221 out220 out219 out218 out217 out216 out215 out214 out213 out212 out211 out210 out209 out208 out207 out206 out205 out204 out203 out202 out201 out200 out199 out198 out197 out196 out195 out194 out193 out192 out191 out190 out189 out188 out187 out186 out185 out184 out183 out182 out181 out180 out179 out178 out177 out176 out175 out174 out173 out172 out171 out170 out169 out168 out167 out166 out165 out164 out163 out162 out161 out160 out159 out158 out157 out156 out155 out154 out153 out152 out151 out150 out149 out148 out147 out146 out145 out144 out143 out142 out141 out140 out139 out138 out137 out136 out135 out134 out133 out132 out131 out130 out129 out128 out127 out126 out125 out124 out123 out122 out121 out120 out119 out118 out117 out116 out115 out114 out113 out112 out111 out110 out109 out108 out107 out106 out105 out104 out103 out102 out101 out100 out99 out98 out97 out96 out95 out94 out93 out92 out91 out90 out89 out88 out87 out86 out85 out84 out83 out82 out81 out80 out79 out78 out77 out76 out75 out74 out73 out72 out71 out70 out69 out68 out67 out66 out65 out64 out63 out62 out61 out60 out59 out58 out57 out56 out55 out54 out53 out52 out51 out50 out49 out48 out47 out46 out45 out44 out43 out42 out41 out40 out39 out38 out37 out36 out35 out34 out33 out32 out31 out30 out29 out28 out27 out26 out25 out24 out23 out22 out21 out20 out19 out18 out17 out16 out15 out14 out13 out12 out11 out10 out9 out8 out7 out6 out5 out4 out3 out2 out1 out0 ldotop_vout ldotop_vdd pass_transistors_256 

.ENDS ldo_core

