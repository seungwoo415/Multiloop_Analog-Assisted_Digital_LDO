
.SUBCKT pass_transistors vg0 vg1 vg2 vg3 vg4 vg5 vg6 vg7 vg8 vg9 vg10 vg11 vg12 vg13 vg14 vg15 vg16 vg17 vg18 vg19 vg20 vg21 vg22 vg23 vg24 vg25 vg26 vg27 vg28 vg29 vg30 vg31 vout vdd 
 
   Xinst1 vout vg0 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst2 vout vg1 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst3 vout vg2 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst4 vout vg3 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst5 vout vg4 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst6 vout vg5 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst7 vout vg6 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst8 vout vg7 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst9 vout vg8 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst10 vout vg9 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst11 vout vg10 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst12 vout vg11 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst13 vout vg12 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst14 vout vg13 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst15 vout vg14 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst16 vout vg15 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst17 vout vg16 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst18 vout vg17 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst19 vout vg18 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst20 vout vg19 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst21 vout vg20 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst22 vout vg21 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst23 vout vg22 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst24 vout vg23 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst25 vout vg24 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst26 vout vg25 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst27 vout vg26 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst28 vout vg27 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst29 vout vg28 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst30 vout vg29 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst31 vout vg30 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst32 vout vg31 vdd vdd sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
.ENDS pass_transistors
