
.SUBCKT pass_transistors Vg_0 Vg_1 Vg_2 Vg_3 Vg_4 Vg_5 Vg_6 Vg_7 Vg_8 Vg_9 Vg_10 Vg_11 Vg_12 Vg_13 Vg_14 Vg_15 Vg_16 Vg_17 Vg_18 Vg_19 Vg_20 Vg_21 Vg_22 Vg_23 Vg_24 Vg_25 Vg_26 Vg_27 Vg_28 Vg_29 Vg_30 Vg_31 Vout VDD 
 
   Xinst1 Vout Vg_0 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst2 Vout Vg_1 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst3 Vout Vg_2 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst4 Vout Vg_3 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst5 Vout Vg_4 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst6 Vout Vg_5 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst7 Vout Vg_6 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst8 Vout Vg_7 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst9 Vout Vg_8 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst10 Vout Vg_9 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst11 Vout Vg_10 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst12 Vout Vg_11 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst13 Vout Vg_12 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst14 Vout Vg_13 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst15 Vout Vg_14 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst16 Vout Vg_15 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst17 Vout Vg_16 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst18 Vout Vg_17 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst19 Vout Vg_18 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst20 Vout Vg_19 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst21 Vout Vg_20 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst22 Vout Vg_21 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst23 Vout Vg_22 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst24 Vout Vg_23 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst25 Vout Vg_24 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst26 Vout Vg_25 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst27 Vout Vg_26 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst28 Vout Vg_27 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst29 Vout Vg_28 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst30 Vout Vg_29 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst31 Vout Vg_30 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
   Xinst32 Vout Vg_31 VDD VDD sky130_fd_pr__pfet_01v8 l=0.25u nf=1 w=1.2u
.ENDS pass_transistors
